
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "pp_loop_interface.svh"
`include "pp_loop_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_TOP.SNR_c_U.if_read;
    assign fifo_intf_1.wr_en = AESL_inst_TOP.SNR_c_U.if_write;
    assign fifo_intf_1.fifo_rd_block = ~(AESL_inst_TOP.AWGN_1_U0.SNR_blk_n);
    assign fifo_intf_1.fifo_wr_block = ~(AESL_inst_TOP.entry_proc_U0.SNR_c_blk_n);
    assign fifo_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_TOP.AES_EN_out_U.if_read;
    assign fifo_intf_2.wr_en = AESL_inst_TOP.AES_EN_out_U.if_write;
    assign fifo_intf_2.fifo_rd_block = ~(AESL_inst_TOP.Modulation_U0.AES_EN_out_blk_n);
    assign fifo_intf_2.fifo_wr_block = ~(AESL_inst_TOP.AES_En_De27_U0.AES_EN_out_blk_n);
    assign fifo_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_TOP.xi_U.if_read;
    assign fifo_intf_3.wr_en = AESL_inst_TOP.xi_U.if_write;
    assign fifo_intf_3.fifo_rd_block = ~(AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.xi_blk_n);
    assign fifo_intf_3.fifo_wr_block = ~(AESL_inst_TOP.Modulation_U0.xi_blk_n);
    assign fifo_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_TOP.xr_U.if_read;
    assign fifo_intf_4.wr_en = AESL_inst_TOP.xr_U.if_write;
    assign fifo_intf_4.fifo_rd_block = ~(AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.xr_blk_n);
    assign fifo_intf_4.fifo_wr_block = ~(AESL_inst_TOP.Modulation_U0.xr_blk_n);
    assign fifo_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_TOP.H_real_U.if_read;
    assign fifo_intf_5.wr_en = AESL_inst_TOP.H_real_U.if_write;
    assign fifo_intf_5.fifo_rd_block = ~(AESL_inst_TOP.split_U0.H_real_blk_n);
    assign fifo_intf_5.fifo_wr_block = ~(AESL_inst_TOP.Rayleigh_1_U0.H_real_blk_n);
    assign fifo_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_TOP.H_imag_U.if_read;
    assign fifo_intf_6.wr_en = AESL_inst_TOP.H_imag_U.if_write;
    assign fifo_intf_6.fifo_rd_block = ~(AESL_inst_TOP.split_1_U0.H_imag_blk_n);
    assign fifo_intf_6.fifo_wr_block = ~(AESL_inst_TOP.Rayleigh_1_U0.H_imag_blk_n);
    assign fifo_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_TOP.H_real_spl0_U.if_read;
    assign fifo_intf_7.wr_en = AESL_inst_TOP.H_real_spl0_U.if_write;
    assign fifo_intf_7.fifo_rd_block = ~(AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.H_real_spl0_blk_n);
    assign fifo_intf_7.fifo_wr_block = ~(AESL_inst_TOP.split_U0.H_real_spl0_blk_n);
    assign fifo_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;
    df_fifo_intf fifo_intf_8(clock,reset);
    assign fifo_intf_8.rd_en = AESL_inst_TOP.H_real_spl1_U.if_read;
    assign fifo_intf_8.wr_en = AESL_inst_TOP.H_real_spl1_U.if_write;
    assign fifo_intf_8.fifo_rd_block = ~(AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.H_real_spl1_blk_n);
    assign fifo_intf_8.fifo_wr_block = ~(AESL_inst_TOP.split_U0.H_real_spl1_blk_n);
    assign fifo_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_8;
    csv_file_dump cstatus_csv_dumper_8;
    df_fifo_monitor fifo_monitor_8;
    df_fifo_intf fifo_intf_9(clock,reset);
    assign fifo_intf_9.rd_en = AESL_inst_TOP.H_imag_spl0_U.if_read;
    assign fifo_intf_9.wr_en = AESL_inst_TOP.H_imag_spl0_U.if_write;
    assign fifo_intf_9.fifo_rd_block = ~(AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.H_imag_spl0_blk_n);
    assign fifo_intf_9.fifo_wr_block = ~(AESL_inst_TOP.split_1_U0.H_imag_spl0_blk_n);
    assign fifo_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_9;
    csv_file_dump cstatus_csv_dumper_9;
    df_fifo_monitor fifo_monitor_9;
    df_fifo_intf fifo_intf_10(clock,reset);
    assign fifo_intf_10.rd_en = AESL_inst_TOP.H_imag_spl1_U.if_read;
    assign fifo_intf_10.wr_en = AESL_inst_TOP.H_imag_spl1_U.if_write;
    assign fifo_intf_10.fifo_rd_block = ~(AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.H_imag_spl1_blk_n);
    assign fifo_intf_10.fifo_wr_block = ~(AESL_inst_TOP.split_1_U0.H_imag_spl1_blk_n);
    assign fifo_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_10;
    csv_file_dump cstatus_csv_dumper_10;
    df_fifo_monitor fifo_monitor_10;
    df_fifo_intf fifo_intf_11(clock,reset);
    assign fifo_intf_11.rd_en = AESL_inst_TOP.R_U.if_read;
    assign fifo_intf_11.wr_en = AESL_inst_TOP.R_U.if_write;
    assign fifo_intf_11.fifo_rd_block = ~(AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.R_blk_n);
    assign fifo_intf_11.fifo_wr_block = ~(AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.R_blk_n);
    assign fifo_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_11;
    csv_file_dump cstatus_csv_dumper_11;
    df_fifo_monitor fifo_monitor_11;
    df_fifo_intf fifo_intf_12(clock,reset);
    assign fifo_intf_12.rd_en = AESL_inst_TOP.Q_U.if_read;
    assign fifo_intf_12.wr_en = AESL_inst_TOP.Q_U.if_write;
    assign fifo_intf_12.fifo_rd_block = ~(AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.Q_blk_n);
    assign fifo_intf_12.fifo_wr_block = ~(AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.Q_blk_n);
    assign fifo_intf_12.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_12;
    csv_file_dump cstatus_csv_dumper_12;
    df_fifo_monitor fifo_monitor_12;
    df_fifo_intf fifo_intf_13(clock,reset);
    assign fifo_intf_13.rd_en = AESL_inst_TOP.channel_out_U.if_read;
    assign fifo_intf_13.wr_en = AESL_inst_TOP.channel_out_U.if_write;
    assign fifo_intf_13.fifo_rd_block = ~(AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.channel_out_blk_n);
    assign fifo_intf_13.fifo_wr_block = ~(AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.channel_out_blk_n);
    assign fifo_intf_13.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_13;
    csv_file_dump cstatus_csv_dumper_13;
    df_fifo_monitor fifo_monitor_13;
    df_fifo_intf fifo_intf_14(clock,reset);
    assign fifo_intf_14.rd_en = AESL_inst_TOP.noise_out_U.if_read;
    assign fifo_intf_14.wr_en = AESL_inst_TOP.noise_out_U.if_write;
    assign fifo_intf_14.fifo_rd_block = ~(AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.noise_out_blk_n);
    assign fifo_intf_14.fifo_wr_block = ~(AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.noise_out_blk_n);
    assign fifo_intf_14.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_14;
    csv_file_dump cstatus_csv_dumper_14;
    df_fifo_monitor fifo_monitor_14;
    df_fifo_intf fifo_intf_15(clock,reset);
    assign fifo_intf_15.rd_en = AESL_inst_TOP.MULQ_out_U.if_read;
    assign fifo_intf_15.wr_en = AESL_inst_TOP.MULQ_out_U.if_write;
    assign fifo_intf_15.fifo_rd_block = ~(AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.MULQ_out_blk_n);
    assign fifo_intf_15.fifo_wr_block = ~(AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.MULQ_out_blk_n);
    assign fifo_intf_15.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_15;
    csv_file_dump cstatus_csv_dumper_15;
    df_fifo_monitor fifo_monitor_15;
    df_fifo_intf fifo_intf_16(clock,reset);
    assign fifo_intf_16.rd_en = AESL_inst_TOP.KB_out_U.if_read;
    assign fifo_intf_16.wr_en = AESL_inst_TOP.KB_out_U.if_write;
    assign fifo_intf_16.fifo_rd_block = ~(AESL_inst_TOP.DeModulation_U0.KB_out_blk_n);
    assign fifo_intf_16.fifo_wr_block = ~(AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.KB_out_blk_n);
    assign fifo_intf_16.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_16;
    csv_file_dump cstatus_csv_dumper_16;
    df_fifo_monitor fifo_monitor_16;
    df_fifo_intf fifo_intf_17(clock,reset);
    assign fifo_intf_17.rd_en = AESL_inst_TOP.demod_out_U.if_read;
    assign fifo_intf_17.wr_en = AESL_inst_TOP.demod_out_U.if_write;
    assign fifo_intf_17.fifo_rd_block = ~(AESL_inst_TOP.AES_En_De_128_U0.demod_out_blk_n);
    assign fifo_intf_17.fifo_wr_block = ~(AESL_inst_TOP.DeModulation_U0.demod_out_blk_n);
    assign fifo_intf_17.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_17;
    csv_file_dump cstatus_csv_dumper_17;
    df_fifo_monitor fifo_monitor_17;

    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_TOP.entry_proc_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_TOP.entry_proc_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_TOP.entry_proc_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_TOP.entry_proc_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_TOP.entry_proc_U0.real_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0 | ~AESL_inst_TOP.entry_proc_U0.SNR_c_blk_n;
    assign process_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_TOP.AES_En_De27_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_TOP.AES_En_De27_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_TOP.AES_En_De27_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_TOP.AES_En_De27_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_TOP.AES_En_De27_U0.real_start;
    assign process_intf_2.pin_stall = 1'b0;
    assign process_intf_2.pout_stall = 1'b0 | ~AESL_inst_TOP.AES_En_De27_U0.AES_EN_out_blk_n;
    assign process_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;
    df_process_intf process_intf_3(clock,reset);
    assign process_intf_3.ap_start = AESL_inst_TOP.Modulation_U0.ap_start;
    assign process_intf_3.ap_ready = AESL_inst_TOP.Modulation_U0.ap_ready;
    assign process_intf_3.ap_done = AESL_inst_TOP.Modulation_U0.ap_done;
    assign process_intf_3.ap_continue = AESL_inst_TOP.Modulation_U0.ap_continue;
    assign process_intf_3.real_start = AESL_inst_TOP.Modulation_U0.real_start;
    assign process_intf_3.pin_stall = 1'b0 | ~AESL_inst_TOP.Modulation_U0.AES_EN_out_blk_n;
    assign process_intf_3.pout_stall = 1'b0 | ~AESL_inst_TOP.Modulation_U0.xi_blk_n | ~AESL_inst_TOP.Modulation_U0.xr_blk_n;
    assign process_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_3;
    csv_file_dump pstatus_csv_dumper_3;
    df_process_monitor process_monitor_3;
    df_process_intf process_intf_4(clock,reset);
    assign process_intf_4.ap_start = AESL_inst_TOP.Rayleigh_1_U0.ap_start;
    assign process_intf_4.ap_ready = AESL_inst_TOP.Rayleigh_1_U0.ap_ready;
    assign process_intf_4.ap_done = AESL_inst_TOP.Rayleigh_1_U0.ap_done;
    assign process_intf_4.ap_continue = AESL_inst_TOP.Rayleigh_1_U0.ap_continue;
    assign process_intf_4.real_start = AESL_inst_TOP.Rayleigh_1_U0.real_start;
    assign process_intf_4.pin_stall = 1'b0;
    assign process_intf_4.pout_stall = 1'b0 | ~AESL_inst_TOP.Rayleigh_1_U0.H_real_blk_n | ~AESL_inst_TOP.Rayleigh_1_U0.H_imag_blk_n;
    assign process_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_4;
    csv_file_dump pstatus_csv_dumper_4;
    df_process_monitor process_monitor_4;
    df_process_intf process_intf_5(clock,reset);
    assign process_intf_5.ap_start = AESL_inst_TOP.split_U0.ap_start;
    assign process_intf_5.ap_ready = AESL_inst_TOP.split_U0.ap_ready;
    assign process_intf_5.ap_done = AESL_inst_TOP.split_U0.ap_done;
    assign process_intf_5.ap_continue = AESL_inst_TOP.split_U0.ap_continue;
    assign process_intf_5.real_start = AESL_inst_TOP.split_U0.real_start;
    assign process_intf_5.pin_stall = 1'b0 | ~AESL_inst_TOP.split_U0.H_real_blk_n;
    assign process_intf_5.pout_stall = 1'b0 | ~AESL_inst_TOP.split_U0.H_real_spl0_blk_n | ~AESL_inst_TOP.split_U0.H_real_spl1_blk_n;
    assign process_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_5;
    csv_file_dump pstatus_csv_dumper_5;
    df_process_monitor process_monitor_5;
    df_process_intf process_intf_6(clock,reset);
    assign process_intf_6.ap_start = AESL_inst_TOP.split_1_U0.ap_start;
    assign process_intf_6.ap_ready = AESL_inst_TOP.split_1_U0.ap_ready;
    assign process_intf_6.ap_done = AESL_inst_TOP.split_1_U0.ap_done;
    assign process_intf_6.ap_continue = AESL_inst_TOP.split_1_U0.ap_continue;
    assign process_intf_6.real_start = AESL_inst_TOP.split_1_U0.ap_start;
    assign process_intf_6.pin_stall = 1'b0 | ~AESL_inst_TOP.split_1_U0.H_imag_blk_n;
    assign process_intf_6.pout_stall = 1'b0 | ~AESL_inst_TOP.split_1_U0.H_imag_spl0_blk_n | ~AESL_inst_TOP.split_1_U0.H_imag_spl1_blk_n;
    assign process_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_6;
    csv_file_dump pstatus_csv_dumper_6;
    df_process_monitor process_monitor_6;
    df_process_intf process_intf_7(clock,reset);
    assign process_intf_7.ap_start = AESL_inst_TOP.QRD_U0.ap_start;
    assign process_intf_7.ap_ready = AESL_inst_TOP.QRD_U0.ap_ready;
    assign process_intf_7.ap_done = AESL_inst_TOP.QRD_U0.ap_done;
    assign process_intf_7.ap_continue = AESL_inst_TOP.QRD_U0.ap_continue;
    assign process_intf_7.real_start = AESL_inst_TOP.QRD_U0.real_start;
    assign process_intf_7.pin_stall = 1'b0 | ~AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.H_real_spl1_blk_n | ~AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.H_imag_spl1_blk_n;
    assign process_intf_7.pout_stall = 1'b0 | ~AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.R_blk_n | ~AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.Q_blk_n;
    assign process_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_7;
    csv_file_dump pstatus_csv_dumper_7;
    df_process_monitor process_monitor_7;
    df_process_intf process_intf_8(clock,reset);
    assign process_intf_8.ap_start = AESL_inst_TOP.channel_mult_U0.ap_start;
    assign process_intf_8.ap_ready = AESL_inst_TOP.channel_mult_U0.ap_ready;
    assign process_intf_8.ap_done = AESL_inst_TOP.channel_mult_U0.ap_done;
    assign process_intf_8.ap_continue = AESL_inst_TOP.channel_mult_U0.ap_continue;
    assign process_intf_8.real_start = AESL_inst_TOP.channel_mult_U0.ap_start;
    assign process_intf_8.pin_stall = 1'b0 | ~AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.H_real_spl0_blk_n | ~AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.H_imag_spl0_blk_n | ~AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.xr_blk_n | ~AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.xi_blk_n;
    assign process_intf_8.pout_stall = 1'b0 | ~AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.channel_out_blk_n;
    assign process_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_8;
    csv_file_dump pstatus_csv_dumper_8;
    df_process_monitor process_monitor_8;
    df_process_intf process_intf_9(clock,reset);
    assign process_intf_9.ap_start = AESL_inst_TOP.AWGN_1_U0.ap_start;
    assign process_intf_9.ap_ready = AESL_inst_TOP.AWGN_1_U0.ap_ready;
    assign process_intf_9.ap_done = AESL_inst_TOP.AWGN_1_U0.ap_done;
    assign process_intf_9.ap_continue = AESL_inst_TOP.AWGN_1_U0.ap_continue;
    assign process_intf_9.real_start = AESL_inst_TOP.AWGN_1_U0.real_start;
    assign process_intf_9.pin_stall = 1'b0 | ~AESL_inst_TOP.AWGN_1_U0.SNR_blk_n | ~AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.channel_out_blk_n;
    assign process_intf_9.pout_stall = 1'b0 | ~AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.noise_out_blk_n;
    assign process_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_9;
    csv_file_dump pstatus_csv_dumper_9;
    df_process_monitor process_monitor_9;
    df_process_intf process_intf_10(clock,reset);
    assign process_intf_10.ap_start = AESL_inst_TOP.matrix_mult_U0.ap_start;
    assign process_intf_10.ap_ready = AESL_inst_TOP.matrix_mult_U0.ap_ready;
    assign process_intf_10.ap_done = AESL_inst_TOP.matrix_mult_U0.ap_done;
    assign process_intf_10.ap_continue = AESL_inst_TOP.matrix_mult_U0.ap_continue;
    assign process_intf_10.real_start = AESL_inst_TOP.matrix_mult_U0.ap_start;
    assign process_intf_10.pin_stall = 1'b0 | ~AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.Q_blk_n | ~AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.noise_out_blk_n;
    assign process_intf_10.pout_stall = 1'b0 | ~AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.MULQ_out_blk_n;
    assign process_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_10;
    csv_file_dump pstatus_csv_dumper_10;
    df_process_monitor process_monitor_10;
    df_process_intf process_intf_11(clock,reset);
    assign process_intf_11.ap_start = AESL_inst_TOP.KBEST_U0.ap_start;
    assign process_intf_11.ap_ready = AESL_inst_TOP.KBEST_U0.ap_ready;
    assign process_intf_11.ap_done = AESL_inst_TOP.KBEST_U0.ap_done;
    assign process_intf_11.ap_continue = AESL_inst_TOP.KBEST_U0.ap_continue;
    assign process_intf_11.real_start = AESL_inst_TOP.KBEST_U0.real_start;
    assign process_intf_11.pin_stall = 1'b0 | ~AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.R_blk_n | ~AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.MULQ_out_blk_n;
    assign process_intf_11.pout_stall = 1'b0 | ~AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.KB_out_blk_n;
    assign process_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_11;
    csv_file_dump pstatus_csv_dumper_11;
    df_process_monitor process_monitor_11;
    df_process_intf process_intf_12(clock,reset);
    assign process_intf_12.ap_start = AESL_inst_TOP.DeModulation_U0.ap_start;
    assign process_intf_12.ap_ready = AESL_inst_TOP.DeModulation_U0.ap_ready;
    assign process_intf_12.ap_done = AESL_inst_TOP.DeModulation_U0.ap_done;
    assign process_intf_12.ap_continue = AESL_inst_TOP.DeModulation_U0.ap_continue;
    assign process_intf_12.real_start = AESL_inst_TOP.DeModulation_U0.real_start;
    assign process_intf_12.pin_stall = 1'b0 | ~AESL_inst_TOP.DeModulation_U0.KB_out_blk_n;
    assign process_intf_12.pout_stall = 1'b0 | ~AESL_inst_TOP.DeModulation_U0.demod_out_blk_n;
    assign process_intf_12.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_12;
    csv_file_dump pstatus_csv_dumper_12;
    df_process_monitor process_monitor_12;
    df_process_intf process_intf_13(clock,reset);
    assign process_intf_13.ap_start = AESL_inst_TOP.AES_En_De_128_U0.ap_start;
    assign process_intf_13.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.ap_ready;
    assign process_intf_13.ap_done = AESL_inst_TOP.AES_En_De_128_U0.ap_done;
    assign process_intf_13.ap_continue = AESL_inst_TOP.AES_En_De_128_U0.ap_continue;
    assign process_intf_13.real_start = AESL_inst_TOP.AES_En_De_128_U0.ap_start;
    assign process_intf_13.pin_stall = 1'b0 | ~AESL_inst_TOP.AES_En_De_128_U0.demod_out_blk_n;
    assign process_intf_13.pout_stall = 1'b0;
    assign process_intf_13.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_13;
    csv_file_dump pstatus_csv_dumper_13;
    df_process_monitor process_monitor_13;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_TOP.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_TOP.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_TOP.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_convertToIntArray_label0_convertToIntArray_label1_fu_284.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_convertToIntArray_label0_convertToIntArray_label1_fu_284.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_convertToIntArray_label0_convertToIntArray_label1_fu_284.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_addRoundKey_fu_322.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_addRoundKey_fu_322.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_addRoundKey_fu_322.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_aes_return_label12_fu_332.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_aes_return_label12_fu_332.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_aes_return_label12_fu_332.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = 1'b0;
    assign module_intf_9.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_aes_return_label12_fu_332.grp_GFMul_fu_342.ap_ready;
    assign module_intf_9.ap_done = 1'b0;
    assign module_intf_9.ap_continue = 1'b0;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = 1'b0;
    assign module_intf_10.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_aes_return_label12_fu_332.grp_GFMul_fu_349.ap_ready;
    assign module_intf_10.ap_done = 1'b0;
    assign module_intf_10.ap_continue = 1'b0;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = 1'b0;
    assign module_intf_11.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_aes_return_label12_fu_332.grp_GFMul_fu_356.ap_ready;
    assign module_intf_11.ap_done = 1'b0;
    assign module_intf_11.ap_continue = 1'b0;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_aes_return_label12_fu_332.grp_addRoundKey_fu_369.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_aes_return_label12_fu_332.grp_addRoundKey_fu_369.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_aes_return_label12_fu_332.grp_addRoundKey_fu_369.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign module_intf_30.ap_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done;
    assign module_intf_30.ap_continue = 1'b1;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_01_fu_3120.ap_start;
    assign module_intf_31.ap_ready = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_01_fu_3120.ap_ready;
    assign module_intf_31.ap_done = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_01_fu_3120.ap_done;
    assign module_intf_31.ap_continue = 1'b1;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_start;
    assign module_intf_32.ap_ready = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_ready;
    assign module_intf_32.ap_done = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_done;
    assign module_intf_32.ap_continue = 1'b1;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_start;
    assign module_intf_33.ap_ready = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_ready;
    assign module_intf_33.ap_done = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_done;
    assign module_intf_33.ap_continue = 1'b1;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_start;
    assign module_intf_34.ap_ready = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_ready;
    assign module_intf_34.ap_done = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_done;
    assign module_intf_34.ap_continue = 1'b1;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_start;
    assign module_intf_35.ap_ready = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_ready;
    assign module_intf_35.ap_done = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_done;
    assign module_intf_35.ap_continue = 1'b1;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_start;
    assign module_intf_36.ap_ready = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_ready;
    assign module_intf_36.ap_done = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_done;
    assign module_intf_36.ap_continue = 1'b1;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.ap_start;
    assign module_intf_37.ap_ready = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.ap_ready;
    assign module_intf_37.ap_done = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.ap_done;
    assign module_intf_37.ap_continue = 1'b1;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_start;
    assign module_intf_38.ap_ready = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ready;
    assign module_intf_38.ap_done = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_done;
    assign module_intf_38.ap_continue = 1'b1;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_start;
    assign module_intf_39.ap_ready = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_ready;
    assign module_intf_39.ap_done = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_done;
    assign module_intf_39.ap_continue = 1'b1;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_start;
    assign module_intf_40.ap_ready = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_ready;
    assign module_intf_40.ap_done = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_done;
    assign module_intf_40.ap_continue = 1'b1;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_start;
    assign module_intf_41.ap_ready = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_ready;
    assign module_intf_41.ap_done = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_done;
    assign module_intf_41.ap_continue = 1'b1;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_1_fu_840.ap_start;
    assign module_intf_42.ap_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_1_fu_840.ap_ready;
    assign module_intf_42.ap_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_1_fu_840.ap_done;
    assign module_intf_42.ap_continue = 1'b1;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;
    nodf_module_intf module_intf_43(clock,reset);
    assign module_intf_43.ap_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_start;
    assign module_intf_43.ap_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_ready;
    assign module_intf_43.ap_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_done;
    assign module_intf_43.ap_continue = 1'b1;
    assign module_intf_43.finish = finish;
    csv_file_dump mstatus_csv_dumper_43;
    nodf_module_monitor module_monitor_43;
    nodf_module_intf module_intf_44(clock,reset);
    assign module_intf_44.ap_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_start;
    assign module_intf_44.ap_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_ready;
    assign module_intf_44.ap_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_done;
    assign module_intf_44.ap_continue = 1'b1;
    assign module_intf_44.finish = finish;
    csv_file_dump mstatus_csv_dumper_44;
    nodf_module_monitor module_monitor_44;
    nodf_module_intf module_intf_45(clock,reset);
    assign module_intf_45.ap_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_start;
    assign module_intf_45.ap_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_ready;
    assign module_intf_45.ap_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_done;
    assign module_intf_45.ap_continue = 1'b1;
    assign module_intf_45.finish = finish;
    csv_file_dump mstatus_csv_dumper_45;
    nodf_module_monitor module_monitor_45;
    nodf_module_intf module_intf_46(clock,reset);
    assign module_intf_46.ap_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_start;
    assign module_intf_46.ap_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_ready;
    assign module_intf_46.ap_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_done;
    assign module_intf_46.ap_continue = 1'b1;
    assign module_intf_46.finish = finish;
    csv_file_dump mstatus_csv_dumper_46;
    nodf_module_monitor module_monitor_46;
    nodf_module_intf module_intf_47(clock,reset);
    assign module_intf_47.ap_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_start;
    assign module_intf_47.ap_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_ready;
    assign module_intf_47.ap_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_done;
    assign module_intf_47.ap_continue = 1'b1;
    assign module_intf_47.finish = finish;
    csv_file_dump mstatus_csv_dumper_47;
    nodf_module_monitor module_monitor_47;
    nodf_module_intf module_intf_48(clock,reset);
    assign module_intf_48.ap_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_75_8_VITIS_LOOP_76_9_fu_1001.ap_start;
    assign module_intf_48.ap_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_75_8_VITIS_LOOP_76_9_fu_1001.ap_ready;
    assign module_intf_48.ap_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_75_8_VITIS_LOOP_76_9_fu_1001.ap_done;
    assign module_intf_48.ap_continue = 1'b1;
    assign module_intf_48.finish = finish;
    csv_file_dump mstatus_csv_dumper_48;
    nodf_module_monitor module_monitor_48;
    nodf_module_intf module_intf_49(clock,reset);
    assign module_intf_49.ap_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_94_11_fu_1070.ap_start;
    assign module_intf_49.ap_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_94_11_fu_1070.ap_ready;
    assign module_intf_49.ap_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_94_11_fu_1070.ap_done;
    assign module_intf_49.ap_continue = 1'b1;
    assign module_intf_49.finish = finish;
    csv_file_dump mstatus_csv_dumper_49;
    nodf_module_monitor module_monitor_49;
    nodf_module_intf module_intf_50(clock,reset);
    assign module_intf_50.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.ap_start;
    assign module_intf_50.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.ap_ready;
    assign module_intf_50.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.ap_done;
    assign module_intf_50.ap_continue = 1'b1;
    assign module_intf_50.finish = finish;
    csv_file_dump mstatus_csv_dumper_50;
    nodf_module_monitor module_monitor_50;
    nodf_module_intf module_intf_51(clock,reset);
    assign module_intf_51.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_start;
    assign module_intf_51.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ready;
    assign module_intf_51.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_done;
    assign module_intf_51.ap_continue = 1'b1;
    assign module_intf_51.finish = finish;
    csv_file_dump mstatus_csv_dumper_51;
    nodf_module_monitor module_monitor_51;
    nodf_module_intf module_intf_52(clock,reset);
    assign module_intf_52.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_start;
    assign module_intf_52.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ready;
    assign module_intf_52.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_done;
    assign module_intf_52.ap_continue = 1'b1;
    assign module_intf_52.finish = finish;
    csv_file_dump mstatus_csv_dumper_52;
    nodf_module_monitor module_monitor_52;
    nodf_module_intf module_intf_53(clock,reset);
    assign module_intf_53.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.ap_start;
    assign module_intf_53.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.ap_ready;
    assign module_intf_53.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.ap_done;
    assign module_intf_53.ap_continue = 1'b1;
    assign module_intf_53.finish = finish;
    csv_file_dump mstatus_csv_dumper_53;
    nodf_module_monitor module_monitor_53;
    nodf_module_intf module_intf_54(clock,reset);
    assign module_intf_54.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_convertToIntArray_label0_convertToIntArray_label1_fu_287.ap_start;
    assign module_intf_54.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_convertToIntArray_label0_convertToIntArray_label1_fu_287.ap_ready;
    assign module_intf_54.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_convertToIntArray_label0_convertToIntArray_label1_fu_287.ap_done;
    assign module_intf_54.ap_continue = 1'b1;
    assign module_intf_54.finish = finish;
    csv_file_dump mstatus_csv_dumper_54;
    nodf_module_monitor module_monitor_54;
    nodf_module_intf module_intf_55(clock,reset);
    assign module_intf_55.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_addRoundKey_label0_fu_325.ap_start;
    assign module_intf_55.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_addRoundKey_label0_fu_325.ap_ready;
    assign module_intf_55.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_addRoundKey_label0_fu_325.ap_done;
    assign module_intf_55.ap_continue = 1'b1;
    assign module_intf_55.finish = finish;
    csv_file_dump mstatus_csv_dumper_55;
    nodf_module_monitor module_monitor_55;
    nodf_module_intf module_intf_56(clock,reset);
    assign module_intf_56.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.ap_start;
    assign module_intf_56.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.ap_ready;
    assign module_intf_56.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.ap_done;
    assign module_intf_56.ap_continue = 1'b1;
    assign module_intf_56.finish = finish;
    csv_file_dump mstatus_csv_dumper_56;
    nodf_module_monitor module_monitor_56;
    nodf_module_intf module_intf_57(clock,reset);
    assign module_intf_57.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_542.ap_start;
    assign module_intf_57.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_542.ap_ready;
    assign module_intf_57.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_542.ap_done;
    assign module_intf_57.ap_continue = 1'b1;
    assign module_intf_57.finish = finish;
    csv_file_dump mstatus_csv_dumper_57;
    nodf_module_monitor module_monitor_57;
    nodf_module_intf module_intf_58(clock,reset);
    assign module_intf_58.ap_start = 1'b0;
    assign module_intf_58.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_542.grp_GFMul_fu_197.ap_ready;
    assign module_intf_58.ap_done = 1'b0;
    assign module_intf_58.ap_continue = 1'b0;
    assign module_intf_58.finish = finish;
    csv_file_dump mstatus_csv_dumper_58;
    nodf_module_monitor module_monitor_58;
    nodf_module_intf module_intf_59(clock,reset);
    assign module_intf_59.ap_start = 1'b0;
    assign module_intf_59.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_542.grp_GFMul_fu_205.ap_ready;
    assign module_intf_59.ap_done = 1'b0;
    assign module_intf_59.ap_continue = 1'b0;
    assign module_intf_59.finish = finish;
    csv_file_dump mstatus_csv_dumper_59;
    nodf_module_monitor module_monitor_59;
    nodf_module_intf module_intf_60(clock,reset);
    assign module_intf_60.ap_start = 1'b0;
    assign module_intf_60.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_542.grp_GFMul_fu_213.ap_ready;
    assign module_intf_60.ap_done = 1'b0;
    assign module_intf_60.ap_continue = 1'b0;
    assign module_intf_60.finish = finish;
    csv_file_dump mstatus_csv_dumper_60;
    nodf_module_monitor module_monitor_60;
    nodf_module_intf module_intf_61(clock,reset);
    assign module_intf_61.ap_start = 1'b0;
    assign module_intf_61.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_542.grp_GFMul_fu_221.ap_ready;
    assign module_intf_61.ap_done = 1'b0;
    assign module_intf_61.ap_continue = 1'b0;
    assign module_intf_61.finish = finish;
    csv_file_dump mstatus_csv_dumper_61;
    nodf_module_monitor module_monitor_61;
    nodf_module_intf module_intf_62(clock,reset);
    assign module_intf_62.ap_start = 1'b0;
    assign module_intf_62.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_542.grp_GFMul_fu_229.ap_ready;
    assign module_intf_62.ap_done = 1'b0;
    assign module_intf_62.ap_continue = 1'b0;
    assign module_intf_62.finish = finish;
    csv_file_dump mstatus_csv_dumper_62;
    nodf_module_monitor module_monitor_62;
    nodf_module_intf module_intf_63(clock,reset);
    assign module_intf_63.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_548.ap_start;
    assign module_intf_63.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_548.ap_ready;
    assign module_intf_63.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_548.ap_done;
    assign module_intf_63.ap_continue = 1'b1;
    assign module_intf_63.finish = finish;
    csv_file_dump mstatus_csv_dumper_63;
    nodf_module_monitor module_monitor_63;
    nodf_module_intf module_intf_64(clock,reset);
    assign module_intf_64.ap_start = 1'b0;
    assign module_intf_64.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_548.grp_GFMul_fu_197.ap_ready;
    assign module_intf_64.ap_done = 1'b0;
    assign module_intf_64.ap_continue = 1'b0;
    assign module_intf_64.finish = finish;
    csv_file_dump mstatus_csv_dumper_64;
    nodf_module_monitor module_monitor_64;
    nodf_module_intf module_intf_65(clock,reset);
    assign module_intf_65.ap_start = 1'b0;
    assign module_intf_65.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_548.grp_GFMul_fu_205.ap_ready;
    assign module_intf_65.ap_done = 1'b0;
    assign module_intf_65.ap_continue = 1'b0;
    assign module_intf_65.finish = finish;
    csv_file_dump mstatus_csv_dumper_65;
    nodf_module_monitor module_monitor_65;
    nodf_module_intf module_intf_66(clock,reset);
    assign module_intf_66.ap_start = 1'b0;
    assign module_intf_66.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_548.grp_GFMul_fu_213.ap_ready;
    assign module_intf_66.ap_done = 1'b0;
    assign module_intf_66.ap_continue = 1'b0;
    assign module_intf_66.finish = finish;
    csv_file_dump mstatus_csv_dumper_66;
    nodf_module_monitor module_monitor_66;
    nodf_module_intf module_intf_67(clock,reset);
    assign module_intf_67.ap_start = 1'b0;
    assign module_intf_67.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_548.grp_GFMul_fu_221.ap_ready;
    assign module_intf_67.ap_done = 1'b0;
    assign module_intf_67.ap_continue = 1'b0;
    assign module_intf_67.finish = finish;
    csv_file_dump mstatus_csv_dumper_67;
    nodf_module_monitor module_monitor_67;
    nodf_module_intf module_intf_68(clock,reset);
    assign module_intf_68.ap_start = 1'b0;
    assign module_intf_68.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deAes_return_label22_fu_332.grp_deMixColumns_fu_548.grp_GFMul_fu_229.ap_ready;
    assign module_intf_68.ap_done = 1'b0;
    assign module_intf_68.ap_continue = 1'b0;
    assign module_intf_68.finish = finish;
    csv_file_dump mstatus_csv_dumper_68;
    nodf_module_monitor module_monitor_68;
    nodf_module_intf module_intf_69(clock,reset);
    assign module_intf_69.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_start;
    assign module_intf_69.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_ready;
    assign module_intf_69.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_done;
    assign module_intf_69.ap_continue = 1'b1;
    assign module_intf_69.finish = finish;
    csv_file_dump mstatus_csv_dumper_69;
    nodf_module_monitor module_monitor_69;
    nodf_module_intf module_intf_70(clock,reset);
    assign module_intf_70.ap_start = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_addRoundKey_label010_fu_349.ap_start;
    assign module_intf_70.ap_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_addRoundKey_label010_fu_349.ap_ready;
    assign module_intf_70.ap_done = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_addRoundKey_label010_fu_349.ap_done;
    assign module_intf_70.ap_continue = 1'b1;
    assign module_intf_70.finish = finish;
    csv_file_dump mstatus_csv_dumper_70;
    nodf_module_monitor module_monitor_70;

    pp_loop_intf #(5) pp_loop_intf_1(clock,reset);
    assign pp_loop_intf_1.pre_loop_state0 = AESL_inst_TOP.Rayleigh_1_U0.ap_ST_fsm_state2;
    assign pp_loop_intf_1.pre_states_valid = 1'b1;
    assign pp_loop_intf_1.post_loop_state0 = AESL_inst_TOP.Rayleigh_1_U0.ap_ST_fsm_state53;
    assign pp_loop_intf_1.post_states_valid = 1'b1;
    assign pp_loop_intf_1.iter_start_state = AESL_inst_TOP.Rayleigh_1_U0.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_start_enable = AESL_inst_TOP.Rayleigh_1_U0.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_1.iter_start_block = AESL_inst_TOP.Rayleigh_1_U0.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.iter_end_state = AESL_inst_TOP.Rayleigh_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_1.iter_end_enable = AESL_inst_TOP.Rayleigh_1_U0.ap_enable_reg_pp0_iter24;
    assign pp_loop_intf_1.iter_end_block = AESL_inst_TOP.Rayleigh_1_U0.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_1.loop_quit_state = AESL_inst_TOP.Rayleigh_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_1.quit_at_end = 1'b1;
    assign pp_loop_intf_1.cur_state = AESL_inst_TOP.Rayleigh_1_U0.ap_CS_fsm;
    assign pp_loop_intf_1.finish = finish;
    csv_file_dump pp_loop_csv_dumper_1;
    pp_loop_monitor #(5) pp_loop_monitor_1;
    seq_loop_intf#(35) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_TOP.AES_En_De27_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_TOP.AES_En_De27_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_1.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.post_loop_state1 = 35'h0;
    assign seq_loop_intf_1.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_TOP.AES_En_De27_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_TOP.AES_En_De27_U0.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_TOP.AES_En_De27_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_TOP.AES_En_De27_U0.ap_ST_fsm_state19;
    assign seq_loop_intf_1.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.iter_end_state1 = AESL_inst_TOP.AES_En_De27_U0.ap_ST_fsm_state35;
    assign seq_loop_intf_1.iter_end_states_valid[1] = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(35) seq_loop_monitor_1;
    seq_loop_intf#(62) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state14;
    assign seq_loop_intf_2.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.post_loop_state1 = 62'h0;
    assign seq_loop_intf_2.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_TOP.QRD_U0.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state13;
    assign seq_loop_intf_2.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.iter_end_state1 = 62'h0;
    assign seq_loop_intf_2.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(62) seq_loop_monitor_2;
    seq_loop_intf#(62) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state30;
    assign seq_loop_intf_3.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.post_loop_state1 = 62'h0;
    assign seq_loop_intf_3.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state14;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_TOP.QRD_U0.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state14;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state29;
    assign seq_loop_intf_3.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.iter_end_state1 = 62'h0;
    assign seq_loop_intf_3.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(62) seq_loop_monitor_3;
    seq_loop_intf#(62) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state31;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state40;
    assign seq_loop_intf_4.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.post_loop_state1 = 62'h0;
    assign seq_loop_intf_4.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state32;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_TOP.QRD_U0.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state32;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state39;
    assign seq_loop_intf_4.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.iter_end_state1 = 62'h0;
    assign seq_loop_intf_4.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(62) seq_loop_monitor_4;
    seq_loop_intf#(62) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state42;
    assign seq_loop_intf_5.pre_states_valid = 1'b1;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state49;
    assign seq_loop_intf_5.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.post_loop_state1 = 62'h0;
    assign seq_loop_intf_5.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state43;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_TOP.QRD_U0.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state43;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state48;
    assign seq_loop_intf_5.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.iter_end_state1 = 62'h0;
    assign seq_loop_intf_5.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(62) seq_loop_monitor_5;
    seq_loop_intf#(62) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state55;
    assign seq_loop_intf_6.pre_states_valid = 1'b1;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state58;
    assign seq_loop_intf_6.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.post_loop_state1 = 62'h0;
    assign seq_loop_intf_6.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state56;
    assign seq_loop_intf_6.quit_states_valid = 1'b1;
    assign seq_loop_intf_6.cur_state = AESL_inst_TOP.QRD_U0.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state56;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_TOP.QRD_U0.ap_ST_fsm_state57;
    assign seq_loop_intf_6.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.iter_end_state1 = 62'h0;
    assign seq_loop_intf_6.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(62) seq_loop_monitor_6;
    seq_loop_intf#(7) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.ap_ST_fsm_state1;
    assign seq_loop_intf_7.pre_states_valid = 1'b1;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.ap_ST_fsm_state5;
    assign seq_loop_intf_7.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.post_loop_state1 = 7'h0;
    assign seq_loop_intf_7.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.ap_ST_fsm_state2;
    assign seq_loop_intf_7.quit_states_valid = 1'b1;
    assign seq_loop_intf_7.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.ap_ST_fsm_state2;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.ap_ST_fsm_state4;
    assign seq_loop_intf_7.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.iter_end_state1 = 7'h0;
    assign seq_loop_intf_7.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(7) seq_loop_monitor_7;
    seq_loop_intf#(7) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.ap_ST_fsm_state1;
    assign seq_loop_intf_8.pre_states_valid = 1'b1;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.ap_ST_fsm_state5;
    assign seq_loop_intf_8.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.post_loop_state1 = 7'h0;
    assign seq_loop_intf_8.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.ap_ST_fsm_state2;
    assign seq_loop_intf_8.quit_states_valid = 1'b1;
    assign seq_loop_intf_8.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.ap_ST_fsm_state2;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.ap_ST_fsm_state4;
    assign seq_loop_intf_8.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.iter_end_state1 = 7'h0;
    assign seq_loop_intf_8.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.one_state_loop = 1'b0;
    assign seq_loop_intf_8.one_state_block = 1'b0;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(7) seq_loop_monitor_8;
    seq_loop_intf#(7) seq_loop_intf_9(clock,reset);
    assign seq_loop_intf_9.pre_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.ap_ST_fsm_state1;
    assign seq_loop_intf_9.pre_states_valid = 1'b1;
    assign seq_loop_intf_9.post_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.ap_ST_fsm_state5;
    assign seq_loop_intf_9.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.post_loop_state1 = 7'h0;
    assign seq_loop_intf_9.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.quit_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.ap_ST_fsm_state2;
    assign seq_loop_intf_9.quit_states_valid = 1'b1;
    assign seq_loop_intf_9.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.ap_CS_fsm;
    assign seq_loop_intf_9.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.ap_ST_fsm_state2;
    assign seq_loop_intf_9.iter_end_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.ap_ST_fsm_state4;
    assign seq_loop_intf_9.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.iter_end_state1 = 7'h0;
    assign seq_loop_intf_9.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.one_state_loop = 1'b0;
    assign seq_loop_intf_9.one_state_block = 1'b0;
    assign seq_loop_intf_9.finish = finish;
    csv_file_dump seq_loop_csv_dumper_9;
    seq_loop_monitor #(7) seq_loop_monitor_9;
    seq_loop_intf#(7) seq_loop_intf_10(clock,reset);
    assign seq_loop_intf_10.pre_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.ap_ST_fsm_state1;
    assign seq_loop_intf_10.pre_states_valid = 1'b1;
    assign seq_loop_intf_10.post_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.ap_ST_fsm_state5;
    assign seq_loop_intf_10.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.post_loop_state1 = 7'h0;
    assign seq_loop_intf_10.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.quit_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.ap_ST_fsm_state2;
    assign seq_loop_intf_10.quit_states_valid = 1'b1;
    assign seq_loop_intf_10.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.ap_CS_fsm;
    assign seq_loop_intf_10.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.ap_ST_fsm_state2;
    assign seq_loop_intf_10.iter_end_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.ap_ST_fsm_state4;
    assign seq_loop_intf_10.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.iter_end_state1 = 7'h0;
    assign seq_loop_intf_10.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.one_state_loop = 1'b0;
    assign seq_loop_intf_10.one_state_block = 1'b0;
    assign seq_loop_intf_10.finish = finish;
    csv_file_dump seq_loop_csv_dumper_10;
    seq_loop_monitor #(7) seq_loop_monitor_10;
    seq_loop_intf#(7) seq_loop_intf_11(clock,reset);
    assign seq_loop_intf_11.pre_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.ap_ST_fsm_state1;
    assign seq_loop_intf_11.pre_states_valid = 1'b1;
    assign seq_loop_intf_11.post_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.ap_ST_fsm_state5;
    assign seq_loop_intf_11.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.post_loop_state1 = 7'h0;
    assign seq_loop_intf_11.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.quit_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.ap_ST_fsm_state2;
    assign seq_loop_intf_11.quit_states_valid = 1'b1;
    assign seq_loop_intf_11.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.ap_CS_fsm;
    assign seq_loop_intf_11.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.ap_ST_fsm_state2;
    assign seq_loop_intf_11.iter_end_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.ap_ST_fsm_state4;
    assign seq_loop_intf_11.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.iter_end_state1 = 7'h0;
    assign seq_loop_intf_11.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.one_state_loop = 1'b0;
    assign seq_loop_intf_11.one_state_block = 1'b0;
    assign seq_loop_intf_11.finish = finish;
    csv_file_dump seq_loop_csv_dumper_11;
    seq_loop_monitor #(7) seq_loop_monitor_11;
    seq_loop_intf#(7) seq_loop_intf_12(clock,reset);
    assign seq_loop_intf_12.pre_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.ap_ST_fsm_state1;
    assign seq_loop_intf_12.pre_states_valid = 1'b1;
    assign seq_loop_intf_12.post_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.ap_ST_fsm_state5;
    assign seq_loop_intf_12.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.post_loop_state1 = 7'h0;
    assign seq_loop_intf_12.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.quit_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.ap_ST_fsm_state2;
    assign seq_loop_intf_12.quit_states_valid = 1'b1;
    assign seq_loop_intf_12.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.ap_CS_fsm;
    assign seq_loop_intf_12.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.ap_ST_fsm_state2;
    assign seq_loop_intf_12.iter_end_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.ap_ST_fsm_state4;
    assign seq_loop_intf_12.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.iter_end_state1 = 7'h0;
    assign seq_loop_intf_12.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.one_state_loop = 1'b0;
    assign seq_loop_intf_12.one_state_block = 1'b0;
    assign seq_loop_intf_12.finish = finish;
    csv_file_dump seq_loop_csv_dumper_12;
    seq_loop_monitor #(7) seq_loop_monitor_12;
    seq_loop_intf#(7) seq_loop_intf_13(clock,reset);
    assign seq_loop_intf_13.pre_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.ap_ST_fsm_state1;
    assign seq_loop_intf_13.pre_states_valid = 1'b1;
    assign seq_loop_intf_13.post_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.ap_ST_fsm_state5;
    assign seq_loop_intf_13.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.post_loop_state1 = 7'h0;
    assign seq_loop_intf_13.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.quit_loop_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.ap_ST_fsm_state2;
    assign seq_loop_intf_13.quit_states_valid = 1'b1;
    assign seq_loop_intf_13.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.ap_CS_fsm;
    assign seq_loop_intf_13.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.ap_ST_fsm_state2;
    assign seq_loop_intf_13.iter_end_state0 = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.ap_ST_fsm_state4;
    assign seq_loop_intf_13.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.iter_end_state1 = 7'h0;
    assign seq_loop_intf_13.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.one_state_loop = 1'b0;
    assign seq_loop_intf_13.one_state_block = 1'b0;
    assign seq_loop_intf_13.finish = finish;
    csv_file_dump seq_loop_csv_dumper_13;
    seq_loop_monitor #(7) seq_loop_monitor_13;
    seq_loop_intf#(20) seq_loop_intf_14(clock,reset);
    assign seq_loop_intf_14.pre_loop_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state9;
    assign seq_loop_intf_14.pre_states_valid = 1'b1;
    assign seq_loop_intf_14.post_loop_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state16;
    assign seq_loop_intf_14.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.post_loop_state1 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state17;
    assign seq_loop_intf_14.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_14.quit_loop_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state10;
    assign seq_loop_intf_14.quit_states_valid = 1'b1;
    assign seq_loop_intf_14.cur_state = AESL_inst_TOP.KBEST_U0.ap_CS_fsm;
    assign seq_loop_intf_14.iter_start_state = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state10;
    assign seq_loop_intf_14.iter_end_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state15;
    assign seq_loop_intf_14.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.iter_end_state1 = 20'h0;
    assign seq_loop_intf_14.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.one_state_loop = 1'b0;
    assign seq_loop_intf_14.one_state_block = 1'b0;
    assign seq_loop_intf_14.finish = finish;
    csv_file_dump seq_loop_csv_dumper_14;
    seq_loop_monitor #(20) seq_loop_monitor_14;
    seq_loop_intf#(20) seq_loop_intf_15(clock,reset);
    assign seq_loop_intf_15.pre_loop_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state6;
    assign seq_loop_intf_15.pre_states_valid = 1'b1;
    assign seq_loop_intf_15.post_loop_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state20;
    assign seq_loop_intf_15.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.post_loop_state1 = 20'h0;
    assign seq_loop_intf_15.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.quit_loop_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state7;
    assign seq_loop_intf_15.quit_states_valid = 1'b1;
    assign seq_loop_intf_15.cur_state = AESL_inst_TOP.KBEST_U0.ap_CS_fsm;
    assign seq_loop_intf_15.iter_start_state = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state7;
    assign seq_loop_intf_15.iter_end_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state19;
    assign seq_loop_intf_15.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.iter_end_state1 = 20'h0;
    assign seq_loop_intf_15.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.one_state_loop = 1'b0;
    assign seq_loop_intf_15.one_state_block = 1'b0;
    assign seq_loop_intf_15.finish = finish;
    csv_file_dump seq_loop_csv_dumper_15;
    seq_loop_monitor #(20) seq_loop_monitor_15;
    seq_loop_intf#(20) seq_loop_intf_16(clock,reset);
    assign seq_loop_intf_16.pre_loop_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state3;
    assign seq_loop_intf_16.pre_states_valid = 1'b1;
    assign seq_loop_intf_16.post_loop_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_16.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.post_loop_state1 = 20'h0;
    assign seq_loop_intf_16.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.quit_loop_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_16.quit_states_valid = 1'b1;
    assign seq_loop_intf_16.cur_state = AESL_inst_TOP.KBEST_U0.ap_CS_fsm;
    assign seq_loop_intf_16.iter_start_state = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state4;
    assign seq_loop_intf_16.iter_end_state0 = AESL_inst_TOP.KBEST_U0.ap_ST_fsm_state20;
    assign seq_loop_intf_16.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.iter_end_state1 = 20'h0;
    assign seq_loop_intf_16.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.one_state_loop = 1'b0;
    assign seq_loop_intf_16.one_state_block = 1'b0;
    assign seq_loop_intf_16.finish = finish;
    csv_file_dump seq_loop_csv_dumper_16;
    seq_loop_monitor #(20) seq_loop_monitor_16;
    seq_loop_intf#(35) seq_loop_intf_17(clock,reset);
    assign seq_loop_intf_17.pre_loop_state0 = AESL_inst_TOP.AES_En_De_128_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_17.pre_states_valid = 1'b1;
    assign seq_loop_intf_17.post_loop_state0 = AESL_inst_TOP.AES_En_De_128_U0.ap_ST_fsm_state1;
    assign seq_loop_intf_17.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.post_loop_state1 = 35'h0;
    assign seq_loop_intf_17.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.quit_loop_state0 = AESL_inst_TOP.AES_En_De_128_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_17.quit_states_valid = 1'b1;
    assign seq_loop_intf_17.cur_state = AESL_inst_TOP.AES_En_De_128_U0.ap_CS_fsm;
    assign seq_loop_intf_17.iter_start_state = AESL_inst_TOP.AES_En_De_128_U0.ap_ST_fsm_state2;
    assign seq_loop_intf_17.iter_end_state0 = AESL_inst_TOP.AES_En_De_128_U0.ap_ST_fsm_state19;
    assign seq_loop_intf_17.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.iter_end_state1 = AESL_inst_TOP.AES_En_De_128_U0.ap_ST_fsm_state35;
    assign seq_loop_intf_17.iter_end_states_valid[1] = 1'b1;
    assign seq_loop_intf_17.one_state_loop = 1'b0;
    assign seq_loop_intf_17.one_state_block = 1'b0;
    assign seq_loop_intf_17.finish = finish;
    csv_file_dump seq_loop_csv_dumper_17;
    seq_loop_monitor #(35) seq_loop_monitor_17;
    upc_loop_intf#(2) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.loop_start = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b0;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(2) upc_loop_monitor_1;
    upc_loop_intf#(6) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.quit_enable = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.loop_start = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_TOP.AES_En_De27_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b0;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(6) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_3.quit_enable = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_3.loop_start = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_TOP.AES_En_De27_U0.grp_aes_return_fu_643.grp_aes_return_Pipeline_subBytes_label0_subBytes_label7_fu_341.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(4) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_TOP.Modulation_U0.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_TOP.Modulation_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_TOP.Modulation_U0.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_4.quit_state = AESL_inst_TOP.Modulation_U0.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_TOP.Modulation_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_TOP.Modulation_U0.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_TOP.Modulation_U0.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_TOP.Modulation_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_TOP.Modulation_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.quit_enable = AESL_inst_TOP.Modulation_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.loop_start = AESL_inst_TOP.Modulation_U0.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_TOP.Modulation_U0.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_TOP.Modulation_U0.ap_done;
    assign upc_loop_intf_4.loop_continue = AESL_inst_TOP.Modulation_U0.ap_continue;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(4) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.quit_enable = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.loop_start = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_TOP.Rayleigh_1_U0.grp_seedInitialization_fu_452.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_TOP.split_U0.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_TOP.split_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_TOP.split_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_TOP.split_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_TOP.split_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_TOP.split_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_TOP.split_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_TOP.split_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_TOP.split_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_TOP.split_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.loop_start = AESL_inst_TOP.split_U0.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_TOP.split_U0.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_TOP.split_U0.ap_done;
    assign upc_loop_intf_6.loop_continue = AESL_inst_TOP.split_U0.ap_continue;
    assign upc_loop_intf_6.quit_at_end = 1'b0;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_TOP.split_1_U0.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_TOP.split_1_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_TOP.split_1_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_TOP.split_1_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_TOP.split_1_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_TOP.split_1_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_TOP.split_1_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_TOP.split_1_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_TOP.split_1_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.quit_enable = AESL_inst_TOP.split_1_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.loop_start = AESL_inst_TOP.split_1_U0.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_TOP.split_1_U0.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_TOP.split_1_U0.ap_done;
    assign upc_loop_intf_7.loop_continue = AESL_inst_TOP.split_1_U0.ap_continue;
    assign upc_loop_intf_7.quit_at_end = 1'b0;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.quit_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.loop_start = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_CHANNEL2REAL_fu_2983.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b0;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.quit_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.loop_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_V_fu_3039.grp_CORDIC_V_Pipeline_VITIS_LOOP_94_2_fu_179.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.quit_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.loop_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3054.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.quit_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.loop_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3072.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;
    upc_loop_intf#(1) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.quit_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.loop_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3081.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b1;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(1) upc_loop_monitor_12;
    upc_loop_intf#(1) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.quit_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.quit_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.loop_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3090.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b1;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(1) upc_loop_monitor_13;
    upc_loop_intf#(1) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.quit_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.quit_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.loop_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3099.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b1;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(1) upc_loop_monitor_14;
    upc_loop_intf#(1) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.quit_state = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.quit_enable = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.loop_start = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_TOP.QRD_U0.grp_CORDIC_R_fu_3108.grp_CORDIC_R_Pipeline_VITIS_LOOP_32_2_fu_163.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b1;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(1) upc_loop_monitor_15;
    upc_loop_intf#(1) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.quit_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.quit_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.loop_start = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_LOOP_02_VITIS_LOOP_260_6_fu_3215.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b0;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(1) upc_loop_monitor_16;
    upc_loop_intf#(27) upc_loop_intf_17(clock,reset);
    assign upc_loop_intf_17.cur_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_CS_fsm;
    assign upc_loop_intf_17.iter_start_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_17.iter_end_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_17.quit_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_17.iter_start_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_17.iter_end_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_17.quit_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_17.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_17.quit_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.loop_start = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_start;
    assign upc_loop_intf_17.loop_ready = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_ready;
    assign upc_loop_intf_17.loop_done = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_277_8_fu_3285.ap_done_int;
    assign upc_loop_intf_17.loop_continue = 1'b1;
    assign upc_loop_intf_17.quit_at_end = 1'b0;
    assign upc_loop_intf_17.finish = finish;
    csv_file_dump upc_loop_csv_dumper_17;
    upc_loop_monitor #(27) upc_loop_monitor_17;
    upc_loop_intf#(1) upc_loop_intf_18(clock,reset);
    assign upc_loop_intf_18.cur_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_CS_fsm;
    assign upc_loop_intf_18.iter_start_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_end_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.quit_state = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_start_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_end_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.quit_block = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_start_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_18.iter_end_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_enable_reg_pp0_iter10;
    assign upc_loop_intf_18.quit_enable = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_enable_reg_pp0_iter10;
    assign upc_loop_intf_18.loop_start = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_start;
    assign upc_loop_intf_18.loop_ready = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_ready;
    assign upc_loop_intf_18.loop_done = AESL_inst_TOP.QRD_U0.grp_QRD_Pipeline_VITIS_LOOP_325_9_VITIS_LOOP_326_10_fu_3420.ap_done_int;
    assign upc_loop_intf_18.loop_continue = 1'b1;
    assign upc_loop_intf_18.quit_at_end = 1'b1;
    assign upc_loop_intf_18.finish = finish;
    csv_file_dump upc_loop_csv_dumper_18;
    upc_loop_monitor #(1) upc_loop_monitor_18;
    upc_loop_intf#(1) upc_loop_intf_19(clock,reset);
    assign upc_loop_intf_19.cur_state = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_CS_fsm;
    assign upc_loop_intf_19.iter_start_state = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_end_state = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.quit_state = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_start_block = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_end_block = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.quit_block = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_start_enable = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.iter_end_enable = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_19.quit_enable = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.loop_start = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_start;
    assign upc_loop_intf_19.loop_ready = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_ready;
    assign upc_loop_intf_19.loop_done = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_CHANNEL2REAL_fu_282.ap_done_int;
    assign upc_loop_intf_19.loop_continue = 1'b1;
    assign upc_loop_intf_19.quit_at_end = 1'b0;
    assign upc_loop_intf_19.finish = finish;
    csv_file_dump upc_loop_csv_dumper_19;
    upc_loop_monitor #(1) upc_loop_monitor_19;
    upc_loop_intf#(8) upc_loop_intf_20(clock,reset);
    assign upc_loop_intf_20.cur_state = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_CS_fsm;
    assign upc_loop_intf_20.iter_start_state = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_end_state = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_ST_fsm_pp0_stage3;
    assign upc_loop_intf_20.quit_state = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_ST_fsm_pp0_stage3;
    assign upc_loop_intf_20.iter_start_block = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_end_block = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_block_pp0_stage3_subdone;
    assign upc_loop_intf_20.quit_block = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_block_pp0_stage3_subdone;
    assign upc_loop_intf_20.iter_start_enable = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_20.iter_end_enable = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_20.quit_enable = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_20.loop_start = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_start;
    assign upc_loop_intf_20.loop_ready = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_ready;
    assign upc_loop_intf_20.loop_done = AESL_inst_TOP.channel_mult_U0.grp_channel_mult_Pipeline_VITIS_LOOP_63_1_fu_354.ap_done_int;
    assign upc_loop_intf_20.loop_continue = 1'b1;
    assign upc_loop_intf_20.quit_at_end = 1'b1;
    assign upc_loop_intf_20.finish = finish;
    csv_file_dump upc_loop_csv_dumper_20;
    upc_loop_monitor #(8) upc_loop_monitor_20;
    upc_loop_intf#(1) upc_loop_intf_21(clock,reset);
    assign upc_loop_intf_21.cur_state = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_CS_fsm;
    assign upc_loop_intf_21.iter_start_state = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_end_state = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.quit_state = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_start_block = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_end_block = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.quit_block = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_start_enable = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_21.iter_end_enable = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_21.quit_enable = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_21.loop_start = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_start;
    assign upc_loop_intf_21.loop_ready = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_ready;
    assign upc_loop_intf_21.loop_done = AESL_inst_TOP.AWGN_1_U0.grp_seedInitialization_fu_58.grp_seedInitialization_Pipeline_SEED_INIT_LOOP_fu_94.ap_done_int;
    assign upc_loop_intf_21.loop_continue = 1'b1;
    assign upc_loop_intf_21.quit_at_end = 1'b1;
    assign upc_loop_intf_21.finish = finish;
    csv_file_dump upc_loop_csv_dumper_21;
    upc_loop_monitor #(1) upc_loop_monitor_21;
    upc_loop_intf#(1) upc_loop_intf_22(clock,reset);
    assign upc_loop_intf_22.cur_state = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_CS_fsm;
    assign upc_loop_intf_22.iter_start_state = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_end_state = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.quit_state = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_start_block = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_end_block = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.quit_block = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_start_enable = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_22.iter_end_enable = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_enable_reg_pp0_iter49;
    assign upc_loop_intf_22.quit_enable = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_enable_reg_pp0_iter49;
    assign upc_loop_intf_22.loop_start = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_start;
    assign upc_loop_intf_22.loop_ready = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_ready;
    assign upc_loop_intf_22.loop_done = AESL_inst_TOP.AWGN_1_U0.grp_AWGN_1_Pipeline_VITIS_LOOP_15_1_fu_72.ap_done_int;
    assign upc_loop_intf_22.loop_continue = 1'b1;
    assign upc_loop_intf_22.quit_at_end = 1'b1;
    assign upc_loop_intf_22.finish = finish;
    csv_file_dump upc_loop_csv_dumper_22;
    upc_loop_monitor #(1) upc_loop_monitor_22;
    upc_loop_intf#(1) upc_loop_intf_23(clock,reset);
    assign upc_loop_intf_23.cur_state = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_CS_fsm;
    assign upc_loop_intf_23.iter_start_state = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_end_state = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.quit_state = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_start_block = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_end_block = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.quit_block = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_start_enable = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_23.iter_end_enable = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_23.quit_enable = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_23.loop_start = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_start;
    assign upc_loop_intf_23.loop_ready = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_ready;
    assign upc_loop_intf_23.loop_done = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_88_1_fu_26.ap_done_int;
    assign upc_loop_intf_23.loop_continue = 1'b1;
    assign upc_loop_intf_23.quit_at_end = 1'b0;
    assign upc_loop_intf_23.finish = finish;
    csv_file_dump upc_loop_csv_dumper_23;
    upc_loop_monitor #(1) upc_loop_monitor_23;
    upc_loop_intf#(8) upc_loop_intf_24(clock,reset);
    assign upc_loop_intf_24.cur_state = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_CS_fsm;
    assign upc_loop_intf_24.iter_start_state = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.iter_end_state = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_ST_fsm_pp0_stage4;
    assign upc_loop_intf_24.quit_state = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_ST_fsm_pp0_stage4;
    assign upc_loop_intf_24.iter_start_block = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.iter_end_block = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_block_pp0_stage4_subdone;
    assign upc_loop_intf_24.quit_block = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_block_pp0_stage4_subdone;
    assign upc_loop_intf_24.iter_start_enable = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_24.iter_end_enable = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_24.quit_enable = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_24.loop_start = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_start;
    assign upc_loop_intf_24.loop_ready = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_ready;
    assign upc_loop_intf_24.loop_done = AESL_inst_TOP.matrix_mult_U0.grp_matrix_mult_Pipeline_VITIS_LOOP_94_2_fu_34.ap_done_int;
    assign upc_loop_intf_24.loop_continue = 1'b1;
    assign upc_loop_intf_24.quit_at_end = 1'b1;
    assign upc_loop_intf_24.finish = finish;
    csv_file_dump upc_loop_csv_dumper_24;
    upc_loop_monitor #(8) upc_loop_monitor_24;
    upc_loop_intf#(1) upc_loop_intf_25(clock,reset);
    assign upc_loop_intf_25.cur_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_CS_fsm;
    assign upc_loop_intf_25.iter_start_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.iter_end_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.quit_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.iter_start_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.iter_end_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.quit_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.iter_start_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_25.iter_end_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_25.quit_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_25.loop_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_start;
    assign upc_loop_intf_25.loop_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_ready;
    assign upc_loop_intf_25.loop_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_21_1_fu_876.ap_done_int;
    assign upc_loop_intf_25.loop_continue = 1'b1;
    assign upc_loop_intf_25.quit_at_end = 1'b0;
    assign upc_loop_intf_25.finish = finish;
    csv_file_dump upc_loop_csv_dumper_25;
    upc_loop_monitor #(1) upc_loop_monitor_25;
    upc_loop_intf#(1) upc_loop_intf_26(clock,reset);
    assign upc_loop_intf_26.cur_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_CS_fsm;
    assign upc_loop_intf_26.iter_start_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.iter_end_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.quit_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.iter_start_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.iter_end_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.quit_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.iter_start_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_26.iter_end_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_26.quit_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_enable_reg_pp0_iter4;
    assign upc_loop_intf_26.loop_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_start;
    assign upc_loop_intf_26.loop_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_ready;
    assign upc_loop_intf_26.loop_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_31_3_fu_884.ap_done_int;
    assign upc_loop_intf_26.loop_continue = 1'b1;
    assign upc_loop_intf_26.quit_at_end = 1'b1;
    assign upc_loop_intf_26.finish = finish;
    csv_file_dump upc_loop_csv_dumper_26;
    upc_loop_monitor #(1) upc_loop_monitor_26;
    upc_loop_intf#(1) upc_loop_intf_27(clock,reset);
    assign upc_loop_intf_27.cur_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_CS_fsm;
    assign upc_loop_intf_27.iter_start_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.iter_end_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.quit_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.iter_start_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.iter_end_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.quit_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.iter_start_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_27.iter_end_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_27.quit_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_27.loop_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_start;
    assign upc_loop_intf_27.loop_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_ready;
    assign upc_loop_intf_27.loop_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_48_5_fu_891.ap_done_int;
    assign upc_loop_intf_27.loop_continue = 1'b1;
    assign upc_loop_intf_27.quit_at_end = 1'b0;
    assign upc_loop_intf_27.finish = finish;
    csv_file_dump upc_loop_csv_dumper_27;
    upc_loop_monitor #(1) upc_loop_monitor_27;
    upc_loop_intf#(1) upc_loop_intf_28(clock,reset);
    assign upc_loop_intf_28.cur_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_CS_fsm;
    assign upc_loop_intf_28.iter_start_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.iter_end_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.quit_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.iter_start_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.iter_end_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.quit_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.iter_start_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_28.iter_end_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_28.quit_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_28.loop_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_start;
    assign upc_loop_intf_28.loop_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_ready;
    assign upc_loop_intf_28.loop_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_104_12_fu_953.ap_done_int;
    assign upc_loop_intf_28.loop_continue = 1'b1;
    assign upc_loop_intf_28.quit_at_end = 1'b0;
    assign upc_loop_intf_28.finish = finish;
    csv_file_dump upc_loop_csv_dumper_28;
    upc_loop_monitor #(1) upc_loop_monitor_28;
    upc_loop_intf#(1) upc_loop_intf_29(clock,reset);
    assign upc_loop_intf_29.cur_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_CS_fsm;
    assign upc_loop_intf_29.iter_start_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.iter_end_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.quit_state = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.iter_start_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.iter_end_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.quit_block = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.iter_start_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_29.iter_end_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_29.quit_enable = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_29.loop_start = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_start;
    assign upc_loop_intf_29.loop_ready = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_ready;
    assign upc_loop_intf_29.loop_done = AESL_inst_TOP.KBEST_U0.grp_KBEST_Pipeline_VITIS_LOOP_57_7_fu_960.ap_done_int;
    assign upc_loop_intf_29.loop_continue = 1'b1;
    assign upc_loop_intf_29.quit_at_end = 1'b0;
    assign upc_loop_intf_29.finish = finish;
    csv_file_dump upc_loop_csv_dumper_29;
    upc_loop_monitor #(1) upc_loop_monitor_29;
    upc_loop_intf#(8) upc_loop_intf_30(clock,reset);
    assign upc_loop_intf_30.cur_state = AESL_inst_TOP.DeModulation_U0.ap_CS_fsm;
    assign upc_loop_intf_30.iter_start_state = AESL_inst_TOP.DeModulation_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.iter_end_state = AESL_inst_TOP.DeModulation_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.quit_state = AESL_inst_TOP.DeModulation_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.iter_start_block = AESL_inst_TOP.DeModulation_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.iter_end_block = AESL_inst_TOP.DeModulation_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.quit_block = AESL_inst_TOP.DeModulation_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.iter_start_enable = AESL_inst_TOP.DeModulation_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_30.iter_end_enable = AESL_inst_TOP.DeModulation_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_30.quit_enable = AESL_inst_TOP.DeModulation_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_30.loop_start = AESL_inst_TOP.DeModulation_U0.ap_start;
    assign upc_loop_intf_30.loop_ready = AESL_inst_TOP.DeModulation_U0.ap_ready;
    assign upc_loop_intf_30.loop_done = AESL_inst_TOP.DeModulation_U0.ap_done;
    assign upc_loop_intf_30.loop_continue = AESL_inst_TOP.DeModulation_U0.ap_continue;
    assign upc_loop_intf_30.quit_at_end = 1'b0;
    assign upc_loop_intf_30.finish = finish;
    csv_file_dump upc_loop_csv_dumper_30;
    upc_loop_monitor #(8) upc_loop_monitor_30;
    upc_loop_intf#(2) upc_loop_intf_31(clock,reset);
    assign upc_loop_intf_31.cur_state = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_CS_fsm;
    assign upc_loop_intf_31.iter_start_state = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.iter_end_state = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.quit_state = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.iter_start_block = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.iter_end_block = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.quit_block = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.iter_start_enable = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_31.iter_end_enable = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_31.quit_enable = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_31.loop_start = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_start;
    assign upc_loop_intf_31.loop_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_ready;
    assign upc_loop_intf_31.loop_done = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label5_fu_12.ap_done_int;
    assign upc_loop_intf_31.loop_continue = 1'b1;
    assign upc_loop_intf_31.quit_at_end = 1'b0;
    assign upc_loop_intf_31.finish = finish;
    csv_file_dump upc_loop_csv_dumper_31;
    upc_loop_monitor #(2) upc_loop_monitor_31;
    upc_loop_intf#(6) upc_loop_intf_32(clock,reset);
    assign upc_loop_intf_32.cur_state = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_CS_fsm;
    assign upc_loop_intf_32.iter_start_state = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_32.iter_end_state = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_32.quit_state = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_32.iter_start_block = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_32.iter_end_block = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_32.quit_block = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_32.iter_start_enable = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_32.iter_end_enable = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_32.quit_enable = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_32.loop_start = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_start;
    assign upc_loop_intf_32.loop_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_ready;
    assign upc_loop_intf_32.loop_done = AESL_inst_TOP.AES_En_De_128_U0.grp_extendKey_fu_633.grp_extendKey_Pipeline_extendKey_label0_fu_20.ap_done_int;
    assign upc_loop_intf_32.loop_continue = 1'b1;
    assign upc_loop_intf_32.quit_at_end = 1'b0;
    assign upc_loop_intf_32.finish = finish;
    csv_file_dump upc_loop_csv_dumper_32;
    upc_loop_monitor #(6) upc_loop_monitor_32;
    upc_loop_intf#(1) upc_loop_intf_33(clock,reset);
    assign upc_loop_intf_33.cur_state = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_CS_fsm;
    assign upc_loop_intf_33.iter_start_state = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.iter_end_state = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.quit_state = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.iter_start_block = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.iter_end_block = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.quit_block = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.iter_start_enable = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_33.iter_end_enable = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_33.quit_enable = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_33.loop_start = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_start;
    assign upc_loop_intf_33.loop_ready = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_ready;
    assign upc_loop_intf_33.loop_done = AESL_inst_TOP.AES_En_De_128_U0.grp_deAes_return_fu_643.grp_deAes_return_Pipeline_deSubBytes_label1_deSubBytes_label13_fu_342.ap_done_int;
    assign upc_loop_intf_33.loop_continue = 1'b1;
    assign upc_loop_intf_33.quit_at_end = 1'b1;
    assign upc_loop_intf_33.finish = finish;
    csv_file_dump upc_loop_csv_dumper_33;
    upc_loop_monitor #(1) upc_loop_monitor_33;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);
    fifo_csv_dumper_8 = new("./depth8.csv");
    cstatus_csv_dumper_8 = new("./chan_status8.csv");
    fifo_monitor_8 = new(fifo_csv_dumper_8,fifo_intf_8,cstatus_csv_dumper_8);
    fifo_csv_dumper_9 = new("./depth9.csv");
    cstatus_csv_dumper_9 = new("./chan_status9.csv");
    fifo_monitor_9 = new(fifo_csv_dumper_9,fifo_intf_9,cstatus_csv_dumper_9);
    fifo_csv_dumper_10 = new("./depth10.csv");
    cstatus_csv_dumper_10 = new("./chan_status10.csv");
    fifo_monitor_10 = new(fifo_csv_dumper_10,fifo_intf_10,cstatus_csv_dumper_10);
    fifo_csv_dumper_11 = new("./depth11.csv");
    cstatus_csv_dumper_11 = new("./chan_status11.csv");
    fifo_monitor_11 = new(fifo_csv_dumper_11,fifo_intf_11,cstatus_csv_dumper_11);
    fifo_csv_dumper_12 = new("./depth12.csv");
    cstatus_csv_dumper_12 = new("./chan_status12.csv");
    fifo_monitor_12 = new(fifo_csv_dumper_12,fifo_intf_12,cstatus_csv_dumper_12);
    fifo_csv_dumper_13 = new("./depth13.csv");
    cstatus_csv_dumper_13 = new("./chan_status13.csv");
    fifo_monitor_13 = new(fifo_csv_dumper_13,fifo_intf_13,cstatus_csv_dumper_13);
    fifo_csv_dumper_14 = new("./depth14.csv");
    cstatus_csv_dumper_14 = new("./chan_status14.csv");
    fifo_monitor_14 = new(fifo_csv_dumper_14,fifo_intf_14,cstatus_csv_dumper_14);
    fifo_csv_dumper_15 = new("./depth15.csv");
    cstatus_csv_dumper_15 = new("./chan_status15.csv");
    fifo_monitor_15 = new(fifo_csv_dumper_15,fifo_intf_15,cstatus_csv_dumper_15);
    fifo_csv_dumper_16 = new("./depth16.csv");
    cstatus_csv_dumper_16 = new("./chan_status16.csv");
    fifo_monitor_16 = new(fifo_csv_dumper_16,fifo_intf_16,cstatus_csv_dumper_16);
    fifo_csv_dumper_17 = new("./depth17.csv");
    cstatus_csv_dumper_17 = new("./chan_status17.csv");
    fifo_monitor_17 = new(fifo_csv_dumper_17,fifo_intf_17,cstatus_csv_dumper_17);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);
    pstall_csv_dumper_3 = new("./stalling3.csv");
    pstatus_csv_dumper_3 = new("./status3.csv");
    process_monitor_3 = new(pstall_csv_dumper_3,process_intf_3,pstatus_csv_dumper_3);
    pstall_csv_dumper_4 = new("./stalling4.csv");
    pstatus_csv_dumper_4 = new("./status4.csv");
    process_monitor_4 = new(pstall_csv_dumper_4,process_intf_4,pstatus_csv_dumper_4);
    pstall_csv_dumper_5 = new("./stalling5.csv");
    pstatus_csv_dumper_5 = new("./status5.csv");
    process_monitor_5 = new(pstall_csv_dumper_5,process_intf_5,pstatus_csv_dumper_5);
    pstall_csv_dumper_6 = new("./stalling6.csv");
    pstatus_csv_dumper_6 = new("./status6.csv");
    process_monitor_6 = new(pstall_csv_dumper_6,process_intf_6,pstatus_csv_dumper_6);
    pstall_csv_dumper_7 = new("./stalling7.csv");
    pstatus_csv_dumper_7 = new("./status7.csv");
    process_monitor_7 = new(pstall_csv_dumper_7,process_intf_7,pstatus_csv_dumper_7);
    pstall_csv_dumper_8 = new("./stalling8.csv");
    pstatus_csv_dumper_8 = new("./status8.csv");
    process_monitor_8 = new(pstall_csv_dumper_8,process_intf_8,pstatus_csv_dumper_8);
    pstall_csv_dumper_9 = new("./stalling9.csv");
    pstatus_csv_dumper_9 = new("./status9.csv");
    process_monitor_9 = new(pstall_csv_dumper_9,process_intf_9,pstatus_csv_dumper_9);
    pstall_csv_dumper_10 = new("./stalling10.csv");
    pstatus_csv_dumper_10 = new("./status10.csv");
    process_monitor_10 = new(pstall_csv_dumper_10,process_intf_10,pstatus_csv_dumper_10);
    pstall_csv_dumper_11 = new("./stalling11.csv");
    pstatus_csv_dumper_11 = new("./status11.csv");
    process_monitor_11 = new(pstall_csv_dumper_11,process_intf_11,pstatus_csv_dumper_11);
    pstall_csv_dumper_12 = new("./stalling12.csv");
    pstatus_csv_dumper_12 = new("./status12.csv");
    process_monitor_12 = new(pstall_csv_dumper_12,process_intf_12,pstatus_csv_dumper_12);
    pstall_csv_dumper_13 = new("./stalling13.csv");
    pstatus_csv_dumper_13 = new("./status13.csv");
    process_monitor_13 = new(pstall_csv_dumper_13,process_intf_13,pstatus_csv_dumper_13);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);
    mstatus_csv_dumper_43 = new("./module_status43.csv");
    module_monitor_43 = new(module_intf_43,mstatus_csv_dumper_43);
    mstatus_csv_dumper_44 = new("./module_status44.csv");
    module_monitor_44 = new(module_intf_44,mstatus_csv_dumper_44);
    mstatus_csv_dumper_45 = new("./module_status45.csv");
    module_monitor_45 = new(module_intf_45,mstatus_csv_dumper_45);
    mstatus_csv_dumper_46 = new("./module_status46.csv");
    module_monitor_46 = new(module_intf_46,mstatus_csv_dumper_46);
    mstatus_csv_dumper_47 = new("./module_status47.csv");
    module_monitor_47 = new(module_intf_47,mstatus_csv_dumper_47);
    mstatus_csv_dumper_48 = new("./module_status48.csv");
    module_monitor_48 = new(module_intf_48,mstatus_csv_dumper_48);
    mstatus_csv_dumper_49 = new("./module_status49.csv");
    module_monitor_49 = new(module_intf_49,mstatus_csv_dumper_49);
    mstatus_csv_dumper_50 = new("./module_status50.csv");
    module_monitor_50 = new(module_intf_50,mstatus_csv_dumper_50);
    mstatus_csv_dumper_51 = new("./module_status51.csv");
    module_monitor_51 = new(module_intf_51,mstatus_csv_dumper_51);
    mstatus_csv_dumper_52 = new("./module_status52.csv");
    module_monitor_52 = new(module_intf_52,mstatus_csv_dumper_52);
    mstatus_csv_dumper_53 = new("./module_status53.csv");
    module_monitor_53 = new(module_intf_53,mstatus_csv_dumper_53);
    mstatus_csv_dumper_54 = new("./module_status54.csv");
    module_monitor_54 = new(module_intf_54,mstatus_csv_dumper_54);
    mstatus_csv_dumper_55 = new("./module_status55.csv");
    module_monitor_55 = new(module_intf_55,mstatus_csv_dumper_55);
    mstatus_csv_dumper_56 = new("./module_status56.csv");
    module_monitor_56 = new(module_intf_56,mstatus_csv_dumper_56);
    mstatus_csv_dumper_57 = new("./module_status57.csv");
    module_monitor_57 = new(module_intf_57,mstatus_csv_dumper_57);
    mstatus_csv_dumper_58 = new("./module_status58.csv");
    module_monitor_58 = new(module_intf_58,mstatus_csv_dumper_58);
    mstatus_csv_dumper_59 = new("./module_status59.csv");
    module_monitor_59 = new(module_intf_59,mstatus_csv_dumper_59);
    mstatus_csv_dumper_60 = new("./module_status60.csv");
    module_monitor_60 = new(module_intf_60,mstatus_csv_dumper_60);
    mstatus_csv_dumper_61 = new("./module_status61.csv");
    module_monitor_61 = new(module_intf_61,mstatus_csv_dumper_61);
    mstatus_csv_dumper_62 = new("./module_status62.csv");
    module_monitor_62 = new(module_intf_62,mstatus_csv_dumper_62);
    mstatus_csv_dumper_63 = new("./module_status63.csv");
    module_monitor_63 = new(module_intf_63,mstatus_csv_dumper_63);
    mstatus_csv_dumper_64 = new("./module_status64.csv");
    module_monitor_64 = new(module_intf_64,mstatus_csv_dumper_64);
    mstatus_csv_dumper_65 = new("./module_status65.csv");
    module_monitor_65 = new(module_intf_65,mstatus_csv_dumper_65);
    mstatus_csv_dumper_66 = new("./module_status66.csv");
    module_monitor_66 = new(module_intf_66,mstatus_csv_dumper_66);
    mstatus_csv_dumper_67 = new("./module_status67.csv");
    module_monitor_67 = new(module_intf_67,mstatus_csv_dumper_67);
    mstatus_csv_dumper_68 = new("./module_status68.csv");
    module_monitor_68 = new(module_intf_68,mstatus_csv_dumper_68);
    mstatus_csv_dumper_69 = new("./module_status69.csv");
    module_monitor_69 = new(module_intf_69,mstatus_csv_dumper_69);
    mstatus_csv_dumper_70 = new("./module_status70.csv");
    module_monitor_70 = new(module_intf_70,mstatus_csv_dumper_70);

    pp_loop_csv_dumper_1 = new("./pp_loop_status1.csv");
    pp_loop_monitor_1 = new(pp_loop_intf_1,pp_loop_csv_dumper_1);


    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);
    seq_loop_csv_dumper_9 = new("./seq_loop_status9.csv");
    seq_loop_monitor_9 = new(seq_loop_intf_9,seq_loop_csv_dumper_9);
    seq_loop_csv_dumper_10 = new("./seq_loop_status10.csv");
    seq_loop_monitor_10 = new(seq_loop_intf_10,seq_loop_csv_dumper_10);
    seq_loop_csv_dumper_11 = new("./seq_loop_status11.csv");
    seq_loop_monitor_11 = new(seq_loop_intf_11,seq_loop_csv_dumper_11);
    seq_loop_csv_dumper_12 = new("./seq_loop_status12.csv");
    seq_loop_monitor_12 = new(seq_loop_intf_12,seq_loop_csv_dumper_12);
    seq_loop_csv_dumper_13 = new("./seq_loop_status13.csv");
    seq_loop_monitor_13 = new(seq_loop_intf_13,seq_loop_csv_dumper_13);
    seq_loop_csv_dumper_14 = new("./seq_loop_status14.csv");
    seq_loop_monitor_14 = new(seq_loop_intf_14,seq_loop_csv_dumper_14);
    seq_loop_csv_dumper_15 = new("./seq_loop_status15.csv");
    seq_loop_monitor_15 = new(seq_loop_intf_15,seq_loop_csv_dumper_15);
    seq_loop_csv_dumper_16 = new("./seq_loop_status16.csv");
    seq_loop_monitor_16 = new(seq_loop_intf_16,seq_loop_csv_dumper_16);
    seq_loop_csv_dumper_17 = new("./seq_loop_status17.csv");
    seq_loop_monitor_17 = new(seq_loop_intf_17,seq_loop_csv_dumper_17);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);
    upc_loop_csv_dumper_17 = new("./upc_loop_status17.csv");
    upc_loop_monitor_17 = new(upc_loop_intf_17,upc_loop_csv_dumper_17);
    upc_loop_csv_dumper_18 = new("./upc_loop_status18.csv");
    upc_loop_monitor_18 = new(upc_loop_intf_18,upc_loop_csv_dumper_18);
    upc_loop_csv_dumper_19 = new("./upc_loop_status19.csv");
    upc_loop_monitor_19 = new(upc_loop_intf_19,upc_loop_csv_dumper_19);
    upc_loop_csv_dumper_20 = new("./upc_loop_status20.csv");
    upc_loop_monitor_20 = new(upc_loop_intf_20,upc_loop_csv_dumper_20);
    upc_loop_csv_dumper_21 = new("./upc_loop_status21.csv");
    upc_loop_monitor_21 = new(upc_loop_intf_21,upc_loop_csv_dumper_21);
    upc_loop_csv_dumper_22 = new("./upc_loop_status22.csv");
    upc_loop_monitor_22 = new(upc_loop_intf_22,upc_loop_csv_dumper_22);
    upc_loop_csv_dumper_23 = new("./upc_loop_status23.csv");
    upc_loop_monitor_23 = new(upc_loop_intf_23,upc_loop_csv_dumper_23);
    upc_loop_csv_dumper_24 = new("./upc_loop_status24.csv");
    upc_loop_monitor_24 = new(upc_loop_intf_24,upc_loop_csv_dumper_24);
    upc_loop_csv_dumper_25 = new("./upc_loop_status25.csv");
    upc_loop_monitor_25 = new(upc_loop_intf_25,upc_loop_csv_dumper_25);
    upc_loop_csv_dumper_26 = new("./upc_loop_status26.csv");
    upc_loop_monitor_26 = new(upc_loop_intf_26,upc_loop_csv_dumper_26);
    upc_loop_csv_dumper_27 = new("./upc_loop_status27.csv");
    upc_loop_monitor_27 = new(upc_loop_intf_27,upc_loop_csv_dumper_27);
    upc_loop_csv_dumper_28 = new("./upc_loop_status28.csv");
    upc_loop_monitor_28 = new(upc_loop_intf_28,upc_loop_csv_dumper_28);
    upc_loop_csv_dumper_29 = new("./upc_loop_status29.csv");
    upc_loop_monitor_29 = new(upc_loop_intf_29,upc_loop_csv_dumper_29);
    upc_loop_csv_dumper_30 = new("./upc_loop_status30.csv");
    upc_loop_monitor_30 = new(upc_loop_intf_30,upc_loop_csv_dumper_30);
    upc_loop_csv_dumper_31 = new("./upc_loop_status31.csv");
    upc_loop_monitor_31 = new(upc_loop_intf_31,upc_loop_csv_dumper_31);
    upc_loop_csv_dumper_32 = new("./upc_loop_status32.csv");
    upc_loop_monitor_32 = new(upc_loop_intf_32,upc_loop_csv_dumper_32);
    upc_loop_csv_dumper_33 = new("./upc_loop_status33.csv");
    upc_loop_monitor_33 = new(upc_loop_intf_33,upc_loop_csv_dumper_33);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(fifo_monitor_8);
    sample_manager_inst.add_one_monitor(fifo_monitor_9);
    sample_manager_inst.add_one_monitor(fifo_monitor_10);
    sample_manager_inst.add_one_monitor(fifo_monitor_11);
    sample_manager_inst.add_one_monitor(fifo_monitor_12);
    sample_manager_inst.add_one_monitor(fifo_monitor_13);
    sample_manager_inst.add_one_monitor(fifo_monitor_14);
    sample_manager_inst.add_one_monitor(fifo_monitor_15);
    sample_manager_inst.add_one_monitor(fifo_monitor_16);
    sample_manager_inst.add_one_monitor(fifo_monitor_17);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(process_monitor_3);
    sample_manager_inst.add_one_monitor(process_monitor_4);
    sample_manager_inst.add_one_monitor(process_monitor_5);
    sample_manager_inst.add_one_monitor(process_monitor_6);
    sample_manager_inst.add_one_monitor(process_monitor_7);
    sample_manager_inst.add_one_monitor(process_monitor_8);
    sample_manager_inst.add_one_monitor(process_monitor_9);
    sample_manager_inst.add_one_monitor(process_monitor_10);
    sample_manager_inst.add_one_monitor(process_monitor_11);
    sample_manager_inst.add_one_monitor(process_monitor_12);
    sample_manager_inst.add_one_monitor(process_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(module_monitor_43);
    sample_manager_inst.add_one_monitor(module_monitor_44);
    sample_manager_inst.add_one_monitor(module_monitor_45);
    sample_manager_inst.add_one_monitor(module_monitor_46);
    sample_manager_inst.add_one_monitor(module_monitor_47);
    sample_manager_inst.add_one_monitor(module_monitor_48);
    sample_manager_inst.add_one_monitor(module_monitor_49);
    sample_manager_inst.add_one_monitor(module_monitor_50);
    sample_manager_inst.add_one_monitor(module_monitor_51);
    sample_manager_inst.add_one_monitor(module_monitor_52);
    sample_manager_inst.add_one_monitor(module_monitor_53);
    sample_manager_inst.add_one_monitor(module_monitor_54);
    sample_manager_inst.add_one_monitor(module_monitor_55);
    sample_manager_inst.add_one_monitor(module_monitor_56);
    sample_manager_inst.add_one_monitor(module_monitor_57);
    sample_manager_inst.add_one_monitor(module_monitor_58);
    sample_manager_inst.add_one_monitor(module_monitor_59);
    sample_manager_inst.add_one_monitor(module_monitor_60);
    sample_manager_inst.add_one_monitor(module_monitor_61);
    sample_manager_inst.add_one_monitor(module_monitor_62);
    sample_manager_inst.add_one_monitor(module_monitor_63);
    sample_manager_inst.add_one_monitor(module_monitor_64);
    sample_manager_inst.add_one_monitor(module_monitor_65);
    sample_manager_inst.add_one_monitor(module_monitor_66);
    sample_manager_inst.add_one_monitor(module_monitor_67);
    sample_manager_inst.add_one_monitor(module_monitor_68);
    sample_manager_inst.add_one_monitor(module_monitor_69);
    sample_manager_inst.add_one_monitor(module_monitor_70);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_9);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_10);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_11);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_12);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_13);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_14);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_15);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_16);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_17);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_17);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_18);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_19);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_20);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_21);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_22);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_23);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_24);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_25);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_26);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_27);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_28);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_29);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_30);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_31);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_32);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_33);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1 || deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
